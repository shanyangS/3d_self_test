module double_top (
	
);

top u0 (

);

top u1(

);

endmodule

