module deserializer (
  input wire t_clk,
  input wire rst_n,

  input wire data_in,
    
  output reg[7:0] data_out
)

reg[3:0] match_reg;


endmodule
